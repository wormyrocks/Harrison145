.title Harrison 145 Main

***** MODELS ***** 
.INCLUDE lib/1812LS.lib
.INCLUDE lib/1812FS.lib
.MODEL MMBT3906 pnp IS=6.84896E-14 BF=135.6 NF=1 BR=0.304 NR=1.0 ISE=5.524807E-13 NE=1.5 ISC=1.71764E-10 NC=1.5 VAF=18.7 VAR=200 IKF=0.0882 IKR=0.229087 RB=1.05 RBM=0.011 IRB=1.51189m RE=0.022 RC=1.57 CJE=8.032025p VJE=0.7118251 MJE=0.3042244 FC=0.5 CJC=9.505229p VJC=0.8414405 MJC=0.5 TF=3.193E-10 ITF=0.4 VTF=4.0 XTF=6 TR=3.342E-8 XTB=1.58 EG=0.78 XTI=3 
.MODEL MMBT3904 NPN IS=4.639f NF=0.9995 ISE=2.091E-14 NE=1.6 BF=160.1 IKF=0.12 VAF=98.69 NR=1.001 ISC=3.257p NC=1.394 BR=5.944 IKR=0.06 VAR=19.29 RB=1 RE=0.3614 RC=1.755 XTB=0 EG=1.11 XTI=3 CJE=5.631p VJE=0.7002 MJE=0.3385 TF=3.001E-10 XTF=27 VTF=1.461 ITF=0.2723 CJC=4.949p VJC=0.5969 MJC=0.1928 XCJC=0.864 TR=9.4E-8 FC=0.5582
.model SM4001 D(Is=14.11n N=1.984 Rs=33.89m Ikf=94.81 Xti=3 Eg=1.11 Cjo=25.89p M=.44 Vj=.3245 Fc=.5 Bv=75 Ibv=10u Tt=5.7u)
.MODEL j2N5484 NJF(Is=.25p Vto=-1.5 Vtotc=-3m Beta=3.0m Lambda=10m Betatce=-.5 Rd=10 Rs=10 Cgs=4p Cgd=4p Kf=3e-17)
.model APot potentiometer( r=10k position=0.5 )
.model d1N914 D(Is=2.52n Rs=.568 N=1.752 Cjo=4p M=.4 tt=20n)
*******************

V1 Vin 0 7.5
V2 V9V 0 9
.include FPO.cir
.include VPO.cir
.include FVO.cir
.include VVO.cir
.include mixer.cir
.include amp.cir 
.include netaliases.cir
.include ctrl.sp
.include display.sp
.end
